//////////////////////////////////////////////////////////////////////////////////
// Company:  Expolog Technologies.
//           Copyright (c) 2023 by Expolog Technologies, Inc. All rights reserved.
//
// Engineer : 
// Revision tag :
// Module Name      :    
// Project Name      : 
// component name : 
// Description: This module provides a test to generate clocks
//              
//
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

//List of Include Files

 `include "cxl_base_test.sv"
`include "req_to_axi_traffic_test.sv"
`include "reset_test.sv"
`include "axi_to_comp_test.sv"
`include "cxlio_FD_test.sv"
`include "cxl_mem_rand_test.sv"
`include "cxl_f2a_rand_test.sv"
