//////////////////////////////////////////////////////////////////////////////////
// Company:  Expolog Technologies.
//           Copyright (c) 2023 by Expolog Technologies, Inc. All rights reserved.
//
// Engineer : 
// Revision tag :
// Module Name      :    
// Project Name      : 
// component name : 
// Description: This module provides a test to generate clocks
//              
//
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
//List of Include Files

  `include "cxl_base_seq.sv"
`include "mem_wr_req.sv"
`include "reset_seq.sv"
`include "axi_to_comp_seq.sv"
`include "req_to_cxlio_FD.sv"
