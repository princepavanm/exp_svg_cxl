//////////////////////////////////////////////////////////////////////////////////
// Company:  Expolog Technologies.
//  Copyright (c) 2023 by Expolog Technologies, Inc. All rights reserved.
//
// Engineer : 
// Revision tag :
// Module Name �: �
// Project Name �: 
// component name : 
// Description: This module provides a test to generate clocks

//
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

class cxl_sbd extends uvm_scoreboard;

  `uvm_analysis_imp_decl(_pcie)

  uvm_analysis_imp_pcie#(pcie_tx, cxl_sbd) imp_pcie_h;

  function new(string name="cxl_sbd", uvm_component parent=null);
    super.new(name, parent);
  endfunction:new

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    imp_pcie_h = new("imp_pcie_h", this);

  endfunction:build_phase

  function void write_pcie(pcie_tx tx);

    `uvm_info("SBD", "Gettting tx from pcie Interface", UVM_LOW)

  endfunction

  virtual task run_phase(uvm_phase phase);
    super.run_phase(phase);

    `uvm_info("SBD","Comparition Logic : Run_phase", UVM_LOW)

  endtask:run_phase

  virtual function check_phase(uvm_phase phase);
    super.check_phase(phase);

    `uvm_info("SBD","Comparition Logic : Check_phase", UVM_LOW)

  endfunction:check_phase

  virtual function report_phase(uvm_phase phase);
    super.report_phase(phase);

    `uvm_info("SBD","Passed and Failed ", UVM_LOW)

  endfunction:report_phase

endclass:cxl_sbd
