//List of Include Files

  `include "cxl_base_test.sv"

