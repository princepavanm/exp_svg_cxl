interface dl_intf(input logic dl_clk, dl_reset_n);

  //Implement Modpot and clocking block here

endinterface:dl_intf
