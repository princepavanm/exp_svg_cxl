interface pass_intf(input logic pass_clk, pass_reset_n);

  //Implement Modpot and clocking block here

endinterface:pass_intf
