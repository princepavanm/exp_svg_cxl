//temp.sv
