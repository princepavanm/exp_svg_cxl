interface arb_intf(input logic arb_clk, arb_reset_n);

  //Implement Modpot and clocking block here

endinterface:arb_intf
