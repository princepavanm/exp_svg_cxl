interface ph_intf(input logic ph_clk, ph_reset_n);

  //Implement Modpot and clocking block here

endinterface:ph_intf
