interface axi_agent_intf(input logic arb_clk, arb_reset_n);

  //Implement Modpot and clocking block here

endinterface:axi_agent_intf
