interface tl_intf(input logic tl_clk, tl_reset_n);

  //Implement Modpot and clocking block here

endinterface:tl_intf
